`define freq    100  // MHz
`define period  1000 / (`freq)  // ns
`define path    "/home/minsu/Desktop/MyVolume/GitLocalRepository/Gitlab/nprc.project/"